// 55:035 sisc processor project
// sisc module

`timescale 1ns/100ps

module sisc (CLK, RST_F, ir);

endmodule
// 55:035 sisc processor project
// test bench for sisc processor

`timescale 1ns/100ps

module sisc_tb;

endmodule
library verilog;
use verilog.vl_types.all;
entity sisc_tb is
end sisc_tb;
